BZh91AY&SY�ë� -*߀Px���������`��������aw��t{���c� 	h.��E���T@�#SDi=h�&eG�ڞ�CM <�G��J��d� @    �&MLL`��J~��6S�i�C�b&�� "Q�)��4��� �h ��D�{Rb2h�� i��!�K�glT�	x -�;�I��fJ��  Y�c,f3&&L�b� R��J��� R�c)fa�z�}���_M��AUЂ�)V~���G(sB�$Q�Q�j㜺]}[j �G�����yeS��1�g3�
�eJ�p 18�EƤ�2<��Ǐ'�x�|�:��<��lN������'Y0u0��%�q��t2O�C�m'��1s�>�O���c]0yn�۬��λu�-��.���үHH���Z�����W�Ħ�^�yW�wmj�[;{�#Yv�.݅�vk���͘����c�,�Mح�n�G)n��[�h�F��.��w�'g��b;w�o"8�,#< ��B� $��#�����&�xF����@��,�[��6�u]$�Z�)�����
2�П��o���7sw�����[os]��������.��vɻԍ���kR7wx���l����V�޷]�1.\���:\�j�$[η�e����o6��0ԛ#Rh�w�N��l���݊�۔���YJ�Lp�sL�D�r��߅�ܨ�g�����M�N
q�܆Hӑ9���I#r )�Jp�rI#�@�q�S�I���@d&8ۑIr�7$����F۞����o�<{��� �Ѫ�-�� �Bk�kj���d10A!0���Q""l�bd�t3��y�#�d	2bS$1�0�J�1+,��m��
F(S1`�H�JR&I��$�LP�1LS��$	 Fٖe����p�$�O8I<�8wnE"od��A6J-&SA��m��F#�sm�s26��H$m2�I�I�Z�Kj��_����j�7�L~ŒN�gé�\Ȅ��̺O:c�r�����x���mӥ��L�0��b�:���f�ڄj��ȴ�d,�F�PQ=��m4��p�	��	��l�Oe�OH��fۍ�v�(�RJ�g�t��hO�Ó��k��9�	�7��pl����ޕ���ݤ��TWL���E����C�Uv^�F��e�����7�DN�UiCwO�O���+��!"`�����*��fe�����������[{��>�E�����<1cA*Ѕ(m#ٓ~�������Ĺw�GW5i��T麂��iӤ���i��3u���Fvc��Xp�I%�4�^<8wP&�M7JfZƕ�DXi�vL4�S��)�ST���)uaãu�&��Pچ����@�x �vg�� Ă�Ą±V��L�#춧��pԏ�����<M>�{"�͹�s��u$���z�Hgy��m�7���7�GR�|�������1a��:n�;�NէN�֑R��a�hV,4����UO7cgN�N��Z�ui��mT�TӇ*֖�;]r�f��;^jci��Ĵ�#Y���L�c��m�<�A�x�}Ti�1����Cni�,Ȏ�ϵ�x��|OV�QI]�"n�E�,�VO;m�"A1������ ���LZ��l�Եfb���w�s �%���$J�ZJ'�A	$��m��I"kkdSȏ�oD$�By$r��hOP�w�܋$a�*�$O9p���A�H����!�m�+�m�s�MNz^"+h�ìyeT��+|r��[1�nI랜�|I;�:5$�[�u���[�ʦ����Lz�܇��=ю�&6���|,���3��p9;gV�NMX�J�]��n'Qݵq���'OR�7�@qw4���\}�D��'
(�b�sHr��n������ 	�?H��n޶���22�[$�Z��e�e���1��[V�l�o��_/d$O���N��G�t���Q9hh��i捕Vrt�]e�Z��{]t4��#4���&"�����Y�m�c��KX��1˶8z�}=i�f�u�yދә/�{��z�ebv��r}����-*X�!9%�a\�eL�G�")"X�k��H�Жs���ňɵ���MA%�"R�ԘT�4:���EO�g<ّ��jXwiy�m!$��Y���{c��a}�h񂁪 � �LE_!�GW`ַ��W��ݗ�)Xn���=Pe}x�b�f��j�v&�~��(�)��x�ӍB��6��|�$-���g�|���2�y��3�,�Cb<�TiD.�^=�#��;SH����|-k>�]dl�<��l��� S
`���"�,EYU"�b���JTc�XAa���Cr���LP�
�{�*eN��n0�A��fï5;��E����j/ 5�T(��_�)�3(�9GyW�v��9�T닗k�l|��$بo(|�;B�>%�5v�$,Mm HL|���V���Z��o��Qͦ����Q����۾bh�\����R��>�xJ�h������ߛ��I"}
i��m�Sf/�L^HiB�āJ��IFn)�Z��J֣WQ���=8ĝ�"
<�G^c��!S����+���ƱYՌۇ�CHă���
8kGk���Q�(���A�����dvUi
�<�ժ���Bޥ�:�ZT]@�v.�ؗA�W��h/�B�ͤ���SQk1B�M: ���	����� "�AChgp��AF�-%�J(��(�Wj�%2��[�L�o�lS��]��BC_�p